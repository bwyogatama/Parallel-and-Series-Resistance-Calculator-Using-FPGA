LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY bcdto7SEG IS
	PORT (bcd : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		HEX: OUT STD_LOGIC_VECTOR (1 TO 7));
END bcdto7SEG;

ARCHITECTURE behavioral OF bcdto7SEG IS

	CONSTANT NOL	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0000";
	CONSTANT SATU	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0001";
	CONSTANT DUA	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0010";
	CONSTANT TIGA	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0011";
	CONSTANT EMPAT	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0100";
	CONSTANT LIMA	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0101";
	CONSTANT ENAM	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0110";
	CONSTANT TUJUH	 : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0111";
	CONSTANT DELAPAN : STD_LOGIC_VECTOR(3 DOWNTO 0)  := "1000";
	CONSTANT SEMBILAN: STD_LOGIC_VECTOR(3 DOWNTO 0)  := "1001";

BEGIN
	
	PROCESS(bcd)
	BEGIN
	CASE bcd IS
	WHEN NOL	=> HEX <="0000001";
	WHEN SATU	=> HEX <="1001111";
	WHEN DUA	=> HEX <="0010010";
	WHEN TIGA	=> HEX <="0000110";
	WHEN EMPAT	=> HEX <="1001100";
	WHEN LIMA	=> HEX <="0100100";
	WHEN ENAM	=> HEX <="0100000";
	WHEN TUJUH	=> HEX <="0001111";
	WHEN DELAPAN	=> HEX <="0000000";
	WHEN SEMBILAN	=> HEX <="0000100";
	WHEN OTHERS	=> HEX <="1111111";
	END CASE;
	END PROCESS;

END behavioral;