LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE components IS

COMPONENT mux2to1
	PORT (w0,w1	:IN STD_LOGIC;
		s		:IN STD_LOGIC;
		f		:OUT STD_LOGIC);
END COMPONENT;


COMPONENT muxdff
			PORT (D0,D1,Sel,Clock 	:IN STD_LOGIC;
					Q					:OUT STD_LOGIC);
END COMPONENT;


COMPONENT regne
	GENERIC(N:INTEGER);
	PORT( 	R		:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
			Resetn	:IN STD_LOGIC;
			E,Clock	:IN STD_LOGIC;
			Q		:OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;
COMPONENT shiftlne
	GENERIC (N:INTEGER);
	PORT (R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0) ;
			L, E, w : IN STD_LOGIC ;
			Clock : IN STD_LOGIC ;
			Q : BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0) ) ;
END COMPONENT ;

COMPONENT shiftrne
	GENERIC ( N : INTEGER  ) ;
	PORT ( R : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0) ;
			L, E, w : IN STD_LOGIC ;
			Clock : IN STD_LOGIC ;
			Q : BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0) ) ;
END COMPONENT ;



COMPONENT downcnt
	GENERIC ( modulus : INTEGER  ) ;
	PORT ( Clock, E, L : IN STD_LOGIC ;
			Q : BUFFER INTEGER RANGE 0 TO modulus-1 ) ;
END COMPONENT ;
COMPONENT bcdto7SEG
	PORT (bcd : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		HEX: OUT STD_LOGIC_VECTOR (1 TO 7));
END COMPONENT;
END components ;